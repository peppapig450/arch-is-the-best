module top;
  initial $display("Arch is the best!");
endmodule
